library verilog;
use verilog.vl_types.all;
entity write_back_stage_sv_unit is
end write_back_stage_sv_unit;
