library verilog;
use verilog.vl_types.all;
entity fetch_stage_sv_unit is
end fetch_stage_sv_unit;
