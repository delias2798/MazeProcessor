library verilog;
use verilog.vl_types.all;
entity memory_stage_sv_unit is
end memory_stage_sv_unit;
