library verilog;
use verilog.vl_types.all;
entity zext_s_sv_unit is
end zext_s_sv_unit;
