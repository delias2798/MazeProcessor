library verilog;
use verilog.vl_types.all;
entity register_control_rom_sv_unit is
end register_control_rom_sv_unit;
