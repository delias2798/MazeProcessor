library verilog;
use verilog.vl_types.all;
entity execute_stage_sv_unit is
end execute_stage_sv_unit;
