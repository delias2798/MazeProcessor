import lc3b_types::*;

module memory_stage
(
	input clk
);

/* Control Signals */

/* Internal Signals */


endmodule: memory_stage