library verilog;
use verilog.vl_types.all;
entity mazeprocessor_sv_unit is
end mazeprocessor_sv_unit;
