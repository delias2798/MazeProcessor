library verilog;
use verilog.vl_types.all;
entity mazeprocessor is
end mazeprocessor;
