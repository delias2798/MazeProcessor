library verilog;
use verilog.vl_types.all;
entity memory_stall_sv_unit is
end memory_stall_sv_unit;
