library verilog;
use verilog.vl_types.all;
entity br_add_sv_unit is
end br_add_sv_unit;
