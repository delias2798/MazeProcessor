library verilog;
use verilog.vl_types.all;
entity decode_stage_sv_unit is
end decode_stage_sv_unit;
