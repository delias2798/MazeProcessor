import lc3b_types::*;

module eviction_wb_datapath
(
	input clk,
	input lc3b_word mem_address,
	input lc3b_data cpu_data,
	input lc3b_data pmem_data,
	input lc3b_word mem_byte_enable,
	
	input valid0_write,
	input valid1_write,
	input valid2_write,
	input valid3_write,
	input valid_in,
	input tag0_write,
	input tag1_write,
	input tag2_write,
	input tag3_write,
	input data0_write,
	input data1_write,
	input data2_write,
	input data3_write,
	input lru_write,
	input [2:0] lru_in,
	input pmem_addr_sig,
	input out_data_sel,
	
	output logic [2:0] lru_out,
	output logic [1:0] cline_and,
	output logic hit,
	output lc3b_data data_out,
	output lc3b_data pdata_out,
	output lc3b_word pmem_address,
	output logic valid0_out,
	output logic valid1_out,
	output logic valid2_out,
	output logic valid3_out
);

lc3b_l2_tag tag;
lc3b_offset offset;

assign tag = mem_address[15:4];
assign offset = mem_address[3:1];

lc3b_l2_tag tag0_out;
lc3b_l2_tag tag1_out;
lc3b_l2_tag tag2_out;
lc3b_l2_tag tag3_out;
lc3b_l2_tag tag_10_out;
lc3b_l2_tag tag_32_out;
lc3b_l2_tag tag_out;
logic comp0_out;
logic comp1_out;
logic comp2_out;
logic comp3_out;

logic cline0_and;
logic cline1_and;
logic cline2_and;
logic cline3_and;

lc3b_data cdata_out;
lc3b_data data0_out;
lc3b_data data1_out;
lc3b_data data2_out;
lc3b_data data3_out;
lc3b_data data_10_out;
lc3b_data data_32_out;

lc3b_word write_back_addr;

/* Valid Arrays */
eviction_wb_array #(.width(1)) valid0
(
	.clk(clk),
	.write(valid0_write),
	.datain(valid_in),
	.dataout(valid0_out)
);

eviction_wb_array #(.width(1)) valid1
(
	.clk(clk),
	.write(valid1_write),
	.datain(valid_in),
	.dataout(valid1_out)
);

eviction_wb_array #(.width(1)) valid2
(
	.clk(clk),
	.write(valid2_write),
	.datain(valid_in),
	.dataout(valid2_out)
);

eviction_wb_array #(.width(1)) valid3
(
	.clk(clk),
	.write(valid3_write),
	.datain(valid_in),
	.dataout(valid3_out)
);

/* LRU Array */
eviction_wb_array #(.width(3)) lru
(
	.clk(clk),
	.write(lru_write),
	.datain(lru_in),
	.dataout(lru_out)
);

/* Tag Arrays */
eviction_wb_array #(.width(8)) tag0
(
	.clk(clk),
	.write(tag0_write),
	.datain(tag),
	.dataout(tag0_out)
);

eviction_wb_array #(.width(8)) tag1
(
	.clk(clk),
	.write(tag1_write),
	.datain(tag),
	.dataout(tag1_out)
);

eviction_wb_array #(.width(8)) tag2
(
	.clk(clk),
	.write(tag2_write),
	.datain(tag),
	.dataout(tag2_out)
);

eviction_wb_array #(.width(8)) tag3
(
	.clk(clk),
	.write(tag3_write),
	.datain(tag),
	.dataout(tag3_out)
);

comparator #(.width(8)) comp0
(
	.value0(tag0_out),
	.value1(tag),
	.out(comp0_out)
);

comparator #(.width(8)) comp1
(
	.value0(tag1_out),
	.value1(tag),
	.out(comp1_out)
);

comparator #(.width(8)) comp2
(
	.value0(tag2_out),
	.value1(tag),
	.out(comp2_out)
);

comparator #(.width(8)) comp3
(
	.value0(tag3_out),
	.value1(tag),
	.out(comp3_out)
);

assign cline0_and = comp0_out & valid0_out;
assign cline1_and = comp1_out & valid1_out;
assign cline2_and = comp2_out & valid2_out;
assign cline3_and = comp3_out & valid3_out;
assign hit = cline0_and | cline1_and | cline2_and | cline3_and;

always_comb
begin
	if (cline0_and)
		cline_and = 2'b00;
	else if (cline1_and)
		cline_and = 2'b01;
	else if (cline2_and)
		cline_and = 2'b10;
	else
		cline_and = 2'b11;
end

eviction_wb_array data0
(
	.clk(clk),
	.write(data0_write),
	.datain(cpu_data),
	.dataout(data0_out)
);

eviction_wb_array data1
(
	.clk(clk),
	.write(data1_write),
	.datain(cpu_data),
	.dataout(data1_out)
);

eviction_wb_array data2
(
	.clk(clk),
	.write(data2_write),
	.datain(cpu_data),
	.dataout(data2_out)
);

eviction_wb_array data3
(
	.clk(clk),
	.write(data3_write),
	.datain(cpu_data),
	.dataout(data3_out)
);

mux4 #(.width(128)) cdata_mux
(
	.sel(cline_and),
	.a(data0_out),
	.b(data1_out),
	.c(data2_out),
	.d(data3_out),
	.f(cdata_out)
);

mux2 #(.width(128)) out_data_mux
(
	.sel(out_data_sel),
	.a(cdata_out),
	.b(pmem_data),
	.f(data_out)
);

/* Address to Physical Memory*/
evict_line evict_data
(
	.a(data0_out),
	.b(data1_out),
	.c(data2_out),
	.d(data3_out),
	.valid_a(valid0_out),
	.valid_b(valid1_out),
	.valid_c(valid2_out),
	.valid_d(valid3_out),
	.lru(lru_out),
	.f(pdata_out)
);

evict_line #(.width(8)) evict_tag
(
	.a(tag0_out),
	.b(tag1_out),
	.c(tag2_out),
	.d(tag3_out),
	.valid_a(valid0_out),
	.valid_b(valid1_out),
	.valid_c(valid2_out),
	.valid_d(valid3_out),
	.lru(lru_out),
	.f(tag_out)
);

assign write_back_addr = {tag_out, 4'b0000};

mux2 #(.width(16)) pmem_addr_mux
(
	.sel(pmem_addr_sig),
	.a(mem_address),
	.b(write_back_addr),
	.f(pmem_address)
);

endmodule: eviction_wb_datapath